/**************************************************************************/
/* code001.v                          For CSC.T341 CLD Archlab TOKYO TECH */
/**************************************************************************/
module main ();
  initial $display("hello, world");
endmodule
