/**************************************************************************/
/* code005.v                          For CSC.T341 CLD Archlab TOKYO TECH */
/**************************************************************************/
/* sample Verilog code */
module main ();
  initial #200 $display("hello, world");
  initial #100 $display("in Verilog HDL");
endmodule
