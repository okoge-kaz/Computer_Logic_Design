/**************************************************************************/
/* code002.v                          For CSC.T341 CLD Archlab TOKYO TECH */
/**************************************************************************/
module main ();
  initial begin
    $display("hello, world");
    $display("in Verilog HDL");
  end
endmodule
