/**************************************************************************/
/* code055.v                          For CSC.T341 CLD Archlab TOKYO TECH */
/**************************************************************************/
`timescale 1ns/100ps
module m_top ();
  reg r_clk=0;
  initial forever #50 r_clk = ~r_clk;
  wire w_out;
  m_main m_main0 (r_clk, w_out);
  initial $dumpfile("main.vcd");
  initial $dumpvars(0, m_main0);
  initial #1000 $finish; 
endmodule


module m_main (w_clk, r_out);
  input  wire w_clk;
  output reg  r_out;

  reg [31:0] r_cnt = 0;
  always@(posedge w_clk) begin
    r_cnt <= (r_cnt==999999) ? 0 : r_cnt +1;
  end

  initial r_out = 0;
  always@(posedge w_clk) begin
    r_out <= (r_cnt==0) ? ~r_out : r_out;
  end
endmodule
