/**************************************************************************/
/* code002_ng.v                       For CSC.T341 CLD Archlab TOKYO TECH */
/**************************************************************************/
module main ();
  initial $display("hello, world");
  $display("in Verilog HDL");
endmodule
